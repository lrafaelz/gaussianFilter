library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity gaussianFilter7x7 is
    port (
        clk     : in std_logic;
        rst     : in std_logic;
        in_0   : in std_logic_vector(15 downto 0);
        in_1   : in std_logic_vector(15 downto 0);
        in_2   : in std_logic_vector(15 downto 0);
        in_3   : in std_logic_vector(15 downto 0);
        in_4   : in std_logic_vector(15 downto 0);
        in_5   : in std_logic_vector(15 downto 0);
        in_6   : in std_logic_vector(15 downto 0);
        in_7   : in std_logic_vector(15 downto 0);
        in_8   : in std_logic_vector(15 downto 0);
        in_9   : in std_logic_vector(15 downto 0);
        in_10   : in std_logic_vector(15 downto 0);
        in_11   : in std_logic_vector(15 downto 0);
        in_12   : in std_logic_vector(15 downto 0);
        in_13   : in std_logic_vector(15 downto 0);
        in_14   : in std_logic_vector(15 downto 0);
        in_15   : in std_logic_vector(15 downto 0);
        in_16   : in std_logic_vector(15 downto 0);
        in_17   : in std_logic_vector(15 downto 0);
        in_18   : in std_logic_vector(15 downto 0);
        in_19   : in std_logic_vector(15 downto 0);
        in_20   : in std_logic_vector(15 downto 0);
        in_21   : in std_logic_vector(15 downto 0);
        in_22   : in std_logic_vector(15 downto 0);
        in_23   : in std_logic_vector(15 downto 0);
        in_24   : in std_logic_vector(15 downto 0);
        in_25   : in std_logic_vector(15 downto 0);
        in_26   : in std_logic_vector(15 downto 0);
        in_27   : in std_logic_vector(15 downto 0);
        in_28   : in std_logic_vector(15 downto 0);
        in_29   : in std_logic_vector(15 downto 0);
        in_30   : in std_logic_vector(15 downto 0);
        in_31   : in std_logic_vector(15 downto 0);
        in_32   : in std_logic_vector(15 downto 0);
        in_33   : in std_logic_vector(15 downto 0);
        in_34   : in std_logic_vector(15 downto 0);
        in_35   : in std_logic_vector(15 downto 0);
        in_36   : in std_logic_vector(15 downto 0);
        in_37   : in std_logic_vector(15 downto 0);
        in_38   : in std_logic_vector(15 downto 0);
        in_39   : in std_logic_vector(15 downto 0);
        in_40   : in std_logic_vector(15 downto 0);
        in_41   : in std_logic_vector(15 downto 0);
        in_42   : in std_logic_vector(15 downto 0);
        in_43   : in std_logic_vector(15 downto 0);
        in_44   : in std_logic_vector(15 downto 0);
        in_45   : in std_logic_vector(15 downto 0);
        in_46   : in std_logic_vector(15 downto 0);
        in_47   : in std_logic_vector(15 downto 0);
        in_48   : in std_logic_vector(15 downto 0);
        out_val : out std_logic_vector(31 downto 0)
        );
        end entity gaussianFilter7x7;
        
        
        architecture behavioral of gaussianFilter7x7 is
            signal out_val_reg          : std_logic_vector(31 downto 0);
            signal partial_product_0    : std_logic_vector(31 downto 0);
            signal partial_product_1    : std_logic_vector(31 downto 0);
            signal partial_product_2    : std_logic_vector(31 downto 0);
            signal partial_product_3    : std_logic_vector(31 downto 0);
            signal partial_product_4    : std_logic_vector(31 downto 0);
            signal partial_product_5    : std_logic_vector(31 downto 0);
            signal partial_product_6    : std_logic_vector(31 downto 0);
            signal partial_product_7    : std_logic_vector(31 downto 0);
            signal partial_product_8    : std_logic_vector(31 downto 0);
            signal partial_product_9    : std_logic_vector(31 downto 0);
            signal partial_product_10   : std_logic_vector(31 downto 0);
            signal partial_product_11   : std_logic_vector(31 downto 0);
            signal partial_product_12   : std_logic_vector(31 downto 0);
            signal partial_product_13   : std_logic_vector(31 downto 0);
            signal partial_product_14   : std_logic_vector(31 downto 0);
            signal partial_product_15   : std_logic_vector(31 downto 0);
            signal partial_product_16   : std_logic_vector(31 downto 0);
            signal partial_product_17   : std_logic_vector(31 downto 0);
            signal partial_product_18   : std_logic_vector(31 downto 0);
            signal partial_product_19   : std_logic_vector(31 downto 0);
            signal partial_product_20   : std_logic_vector(31 downto 0);
            signal partial_product_21   : std_logic_vector(31 downto 0);
            signal partial_product_22   : std_logic_vector(31 downto 0);
            signal partial_product_23   : std_logic_vector(31 downto 0);
            signal partial_product_24   : std_logic_vector(31 downto 0);
            signal partial_product_25   : std_logic_vector(31 downto 0);
            signal partial_product_26   : std_logic_vector(31 downto 0);
            signal partial_product_27   : std_logic_vector(31 downto 0);
            signal partial_product_28   : std_logic_vector(31 downto 0);
            signal partial_product_29   : std_logic_vector(31 downto 0);
            signal partial_product_30   : std_logic_vector(31 downto 0);
            signal partial_product_31   : std_logic_vector(31 downto 0);
            signal partial_product_32   : std_logic_vector(31 downto 0);
            signal partial_product_33   : std_logic_vector(31 downto 0);
            signal partial_product_34   : std_logic_vector(31 downto 0);
            signal partial_product_35   : std_logic_vector(31 downto 0);
            signal partial_product_36   : std_logic_vector(31 downto 0);
            signal partial_product_37   : std_logic_vector(31 downto 0);
            signal partial_product_38   : std_logic_vector(31 downto 0);
            signal partial_product_39   : std_logic_vector(31 downto 0);
            signal partial_product_40   : std_logic_vector(31 downto 0);
            signal partial_product_41   : std_logic_vector(31 downto 0);
            signal partial_product_42   : std_logic_vector(31 downto 0);
            signal partial_product_43   : std_logic_vector(31 downto 0);
            signal partial_product_44   : std_logic_vector(31 downto 0);
            signal partial_product_45   : std_logic_vector(31 downto 0);
            signal partial_product_46   : std_logic_vector(31 downto 0);
            signal partial_product_47   : std_logic_vector(31 downto 0);
            signal partial_product_48   : std_logic_vector(31 downto 0);

            -- input registers
            signal in0_reg              : std_logic_vector(15 downto 0);
            signal in1_reg              : std_logic_vector(15 downto 0);
            signal in2_reg              : std_logic_vector(15 downto 0);
            signal in3_reg              : std_logic_vector(15 downto 0);
            signal in4_reg              : std_logic_vector(15 downto 0);
            signal in5_reg              : std_logic_vector(15 downto 0);
            signal in6_reg              : std_logic_vector(15 downto 0);
            signal in7_reg              : std_logic_vector(15 downto 0);
            signal in8_reg              : std_logic_vector(15 downto 0);
            signal in9_reg              : std_logic_vector(15 downto 0);
            signal in10_reg             : std_logic_vector(15 downto 0);
            signal in11_reg             : std_logic_vector(15 downto 0);
            signal in12_reg             : std_logic_vector(15 downto 0);
            signal in13_reg             : std_logic_vector(15 downto 0);
            signal in14_reg             : std_logic_vector(15 downto 0);
            signal in15_reg             : std_logic_vector(15 downto 0);
            signal in16_reg             : std_logic_vector(15 downto 0);
            signal in17_reg             : std_logic_vector(15 downto 0);
            signal in18_reg             : std_logic_vector(15 downto 0);
            signal in19_reg             : std_logic_vector(15 downto 0);
            signal in20_reg             : std_logic_vector(15 downto 0);
            signal in21_reg             : std_logic_vector(15 downto 0);
            signal in22_reg             : std_logic_vector(15 downto 0);
            signal in23_reg             : std_logic_vector(15 downto 0);
            signal in24_reg             : std_logic_vector(15 downto 0);
            signal in25_reg             : std_logic_vector(15 downto 0);
            signal in26_reg             : std_logic_vector(15 downto 0);
            signal in27_reg             : std_logic_vector(15 downto 0);
            signal in28_reg             : std_logic_vector(15 downto 0);
            signal in29_reg             : std_logic_vector(15 downto 0);
            signal in30_reg             : std_logic_vector(15 downto 0);
            signal in31_reg             : std_logic_vector(15 downto 0);
            signal in32_reg             : std_logic_vector(15 downto 0);
            signal in33_reg             : std_logic_vector(15 downto 0);
            signal in34_reg             : std_logic_vector(15 downto 0);
            signal in35_reg             : std_logic_vector(15 downto 0);
            signal in36_reg             : std_logic_vector(15 downto 0);
            signal in37_reg             : std_logic_vector(15 downto 0);
            signal in38_reg             : std_logic_vector(15 downto 0);
            signal in39_reg             : std_logic_vector(15 downto 0);
            signal in40_reg             : std_logic_vector(15 downto 0);
            signal in41_reg             : std_logic_vector(15 downto 0);
            signal in42_reg             : std_logic_vector(15 downto 0);
            signal in43_reg             : std_logic_vector(15 downto 0);
            signal in44_reg             : std_logic_vector(15 downto 0);
            signal in45_reg             : std_logic_vector(15 downto 0);
            signal in46_reg             : std_logic_vector(15 downto 0);
            signal in47_reg             : std_logic_vector(15 downto 0);
            signal in48_reg             : std_logic_vector(15 downto 0);
            
            begin
            process(clk, rst)
            begin
                if rst = '1' then
                    out_val_reg <= (others => '0');
                    in0_reg <= (others => '0');
                    in1_reg <= (others => '0');
                    in2_reg <= (others => '0');
                    in3_reg <= (others => '0');
                    in4_reg <= (others => '0');
                    in5_reg <= (others => '0');
                    in6_reg <= (others => '0');
                    in7_reg <= (others => '0');
                    in8_reg <= (others => '0');
                    in9_reg <= (others => '0');
                    in10_reg <= (others => '0');
                    in11_reg <= (others => '0');
                    in12_reg <= (others => '0');
                    in13_reg <= (others => '0');
                    in14_reg <= (others => '0');
                    in15_reg <= (others => '0');
                    in16_reg <= (others => '0');
                    in17_reg <= (others => '0');
                    in18_reg <= (others => '0');
                    in19_reg <= (others => '0');
                    in20_reg <= (others => '0');
                    in21_reg <= (others => '0');
                    in22_reg <= (others => '0');
                    in23_reg <= (others => '0');
                    in24_reg <= (others => '0');
                    in25_reg <= (others => '0');
                    in26_reg <= (others => '0');
                    in27_reg <= (others => '0');
                    in28_reg <= (others => '0');
                    in29_reg <= (others => '0');
                    in30_reg <= (others => '0');
                    in31_reg <= (others => '0');
                    in32_reg <= (others => '0');
                    in33_reg <= (others => '0');
                    in34_reg <= (others => '0');
                    in35_reg <= (others => '0');
                    in36_reg <= (others => '0');
                    in37_reg <= (others => '0');
                    in38_reg <= (others => '0');
                    in39_reg <= (others => '0');
                    in40_reg <= (others => '0');
                    in41_reg <= (others => '0');
                    in42_reg <= (others => '0');
                    in43_reg <= (others => '0');
                    in44_reg <= (others => '0');
                    in45_reg <= (others => '0');
                    in46_reg <= (others => '0');
                    in47_reg <= (others => '0');
                    in48_reg <= (others => '0');

                elsif rising_edge(clk) then
                    -- INPUT REGISTERS
                    in0_reg <= in_0;
                    in1_reg <= in_1;
                    in2_reg <= in_2;
                    in3_reg <= in_3;
                    in4_reg <= in_4;
                    in5_reg <= in_5;
                    in6_reg <= in_6;
                    in7_reg <= in_7;
                    in8_reg <= in_8;
                    in9_reg <= in_9;
                    in10_reg <= in_10;
                    in11_reg <= in_11;
                    in12_reg <= in_12;
                    in13_reg <= in_13;
                    in14_reg <= in_14;
                    in15_reg <= in_15;
                    in16_reg <= in_16;
                    in17_reg <= in_17;
                    in18_reg <= in_18;
                    in19_reg <= in_19;
                    in20_reg <= in_20;
                    in21_reg <= in_21;
                    in22_reg <= in_22;
                    in23_reg <= in_23;
                    in24_reg <= in_24;
                    in25_reg <= in_25;
                    in26_reg <= in_26;
                    in27_reg <= in_27;
                    in28_reg <= in_28;
                    in29_reg <= in_29;
                    in30_reg <= in_30;
                    in31_reg <= in_31;
                    in32_reg <= in_32;
                    in33_reg <= in_33;
                    in34_reg <= in_34;
                    in35_reg <= in_35;
                    in36_reg <= in_36;
                    in37_reg <= in_37;
                    in38_reg <= in_38;
                    in39_reg <= in_39;
                    in40_reg <= in_40;
                    in41_reg <= in_41;
                    in42_reg <= in_42;
                    in43_reg <= in_43;
                    in44_reg <= in_44;
                    in45_reg <= in_45;
                    in46_reg <= in_46;
                    in47_reg <= in_47;
                    in48_reg <= in_48;

                    -- SUM
                    out_val_reg <= std_logic_vector(unsigned(partial_product_0) + unsigned(partial_product_1) + unsigned(partial_product_2) + unsigned(partial_product_3) + unsigned(partial_product_4) + unsigned(partial_product_5) + unsigned(partial_product_6) + unsigned(partial_product_7) + unsigned(partial_product_8) + unsigned(partial_product_9) + unsigned(partial_product_10) + unsigned(partial_product_11) + unsigned(partial_product_12) + unsigned(partial_product_13) + unsigned(partial_product_14) + unsigned(partial_product_15) + unsigned(partial_product_16) + unsigned(partial_product_17) + unsigned(partial_product_18) + unsigned(partial_product_19) + unsigned(partial_product_20) + unsigned(partial_product_21) + unsigned(partial_product_22) + unsigned(partial_product_23) + unsigned(partial_product_24) + unsigned(partial_product_25) + unsigned(partial_product_26) + unsigned(partial_product_27) + unsigned(partial_product_28) + unsigned(partial_product_29) + unsigned(partial_product_30) + unsigned(partial_product_31) + unsigned(partial_product_32) + unsigned(partial_product_33) + unsigned(partial_product_34) + unsigned(partial_product_35) + unsigned(partial_product_36) + unsigned(partial_product_37) + unsigned(partial_product_38) + unsigned(partial_product_39) + unsigned(partial_product_40) + unsigned(partial_product_41) + unsigned(partial_product_42) + unsigned(partial_product_43) + unsigned(partial_product_44) + unsigned(partial_product_45) + unsigned(partial_product_46) + unsigned(partial_product_47) + unsigned(partial_product_48));

                end if;
            end process;
            -- (0, 0)
            partial_product_0 <= std_logic_vector(unsigned(in0_reg) * 0);
            partial_product_1 <= std_logic_vector(unsigned(in1_reg) * 1);
            partial_product_2 <= std_logic_vector(unsigned(in2_reg) * 1);
            partial_product_3 <= std_logic_vector(unsigned(in3_reg) * 1);
            partial_product_4 <= std_logic_vector(unsigned(in4_reg) * 1);
            partial_product_5 <= std_logic_vector(unsigned(in5_reg) * 1);
            partial_product_6 <= std_logic_vector(unsigned(in6_reg) * 0);
            -- (1, 0)
            partial_product_7 <= std_logic_vector(unsigned(in7_reg) * 1);
            partial_product_8 <= std_logic_vector(unsigned(in8_reg) * 2);
            partial_product_9 <= std_logic_vector(unsigned(in9_reg) * 4);
            partial_product_10 <= std_logic_vector(unsigned(in10_reg) * 5);
            partial_product_11 <= std_logic_vector(unsigned(in11_reg) * 4);
            partial_product_12 <= std_logic_vector(unsigned(in12_reg) * 2);
            partial_product_13 <= std_logic_vector(unsigned(in13_reg) * 1);
            -- (2, 0)
            partial_product_14 <= std_logic_vector(unsigned(in14_reg) * 1);
            partial_product_15 <= std_logic_vector(unsigned(in15_reg) * 4);
            partial_product_16 <= std_logic_vector(unsigned(in16_reg) * 8);
            partial_product_17 <= std_logic_vector(unsigned(in17_reg) * 10);
            partial_product_18 <= std_logic_vector(unsigned(in18_reg) * 8);
            partial_product_19 <= std_logic_vector(unsigned(in19_reg) * 4);
            partial_product_20 <= std_logic_vector(unsigned(in20_reg) * 1);
            -- (3, 0)
            partial_product_21 <= std_logic_vector(unsigned(in21_reg) * 1);
            partial_product_22 <= std_logic_vector(unsigned(in22_reg) * 5);
            partial_product_23 <= std_logic_vector(unsigned(in23_reg) * 10);
            partial_product_24 <= std_logic_vector(unsigned(in24_reg) * 13);
            partial_product_25 <= std_logic_vector(unsigned(in25_reg) * 10);
            partial_product_26 <= std_logic_vector(unsigned(in26_reg) * 5);
            partial_product_27 <= std_logic_vector(unsigned(in27_reg) * 1);
            -- (4, 0)
            partial_product_28 <= std_logic_vector(unsigned(in28_reg) * 1);
            partial_product_29 <= std_logic_vector(unsigned(in29_reg) * 4);
            partial_product_30 <= std_logic_vector(unsigned(in30_reg) * 8);
            partial_product_31 <= std_logic_vector(unsigned(in31_reg) * 10);
            partial_product_32 <= std_logic_vector(unsigned(in32_reg) * 8);
            partial_product_33 <= std_logic_vector(unsigned(in33_reg) * 4);
            partial_product_34 <= std_logic_vector(unsigned(in34_reg) * 1);
            -- (5, 0)
            partial_product_35 <= std_logic_vector(unsigned(in35_reg) * 1);
            partial_product_36 <= std_logic_vector(unsigned(in36_reg) * 2);
            partial_product_37 <= std_logic_vector(unsigned(in37_reg) * 4);
            partial_product_38 <= std_logic_vector(unsigned(in38_reg) * 5);
            partial_product_39 <= std_logic_vector(unsigned(in39_reg) * 4);
            partial_product_40 <= std_logic_vector(unsigned(in40_reg) * 2);
            partial_product_41 <= std_logic_vector(unsigned(in41_reg) * 1);
            -- (6, 0)
            partial_product_42 <= std_logic_vector(unsigned(in42_reg) * 0);
            partial_product_43 <= std_logic_vector(unsigned(in43_reg) * 1);
            partial_product_44 <= std_logic_vector(unsigned(in44_reg) * 1);
            partial_product_45 <= std_logic_vector(unsigned(in45_reg) * 1);
            partial_product_46 <= std_logic_vector(unsigned(in46_reg) * 1);
            partial_product_47 <= std_logic_vector(unsigned(in47_reg) * 1);
            partial_product_48 <= std_logic_vector(unsigned(in48_reg) * 0);


            out_val <= out_val_reg;
    end architecture behavioral;
    